-- PLL.vhd

-- Generated using ACDS version 13.0sp1 232 at 2017.05.27.21:50:13

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL is
	port (
		clock_27_clk    : in  std_logic := '0'; --    clock_27.clk
		pixel_clock_clk : out std_logic;        -- pixel_clock.clk
		reset_reset     : in  std_logic := '0'  --       reset.reset
	);
end entity PLL;

architecture rtl of PLL is
	component PLL_PLL is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component PLL_PLL;

begin

	pll : component PLL_PLL
		port map (
			clk       => clock_27_clk,    --       inclk_interface.clk
			reset     => reset_reset,     -- inclk_interface_reset.reset
			read      => open,            --             pll_slave.read
			write     => open,            --                      .write
			address   => open,            --                      .address
			readdata  => open,            --                      .readdata
			writedata => open,            --                      .writedata
			c0        => pixel_clock_clk, --                    c0.clk
			areset    => open,            --        areset_conduit.export
			locked    => open,            --        locked_conduit.export
			phasedone => open             --     phasedone_conduit.export
		);

end architecture rtl; -- of PLL
